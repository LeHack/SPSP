package sm410564_formats is
    type data_display_formats is (decimal, mixed, hexadecimal);
end package;
